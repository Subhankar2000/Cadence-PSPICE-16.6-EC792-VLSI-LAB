123_Amrita EXP-1(c) CMOS Two input NAND Gate DT-04112020
vdd 1 0 DC 5v
va 2 0 PULSE 0 5 0 0.1ns 0.1ns 50ns 100ns
vb 3 0 PULSE 0 5 0 0.1ns 0.1ns 100ns 200ns
m1 4 2 1 1 pmod(w=40u l=10u)
m2 4 3 1 1 pmod(w=40u l=10u)
m3 4 2 5 5 nmod(w=10u l=2u)
m4 5 3 0 0 nmod(w=10u l=2u)
.MODEL pmod pmos(vto = -1 lambda=0.02)
.MODEL nmod nmos(vto =  1 lambda=0.02)
.TRAN 0ns 600ns
.PROBE
.END