EXP-1(a) CMOS Inverters with varying Kn(div by)Kp [29-Subhankar Karmakar]A11 DT-04092020
v1 1 0 DC 0
v2 5 0 DC 5
m1 2 1 5 5 pmod(w=10u  l=10u)
m2 3 1 5 5 pmod(w=10u  l=10u)
m3 4 1 5 5 pmod(w=10u  l=10u)
m4 2 1 0 0 nmod(w=200u l=2u)
m5 3 1 0 0 nmod(w=20u  l=2u)
m6 4 1 0 0 nmod(w=2u   l=2u)
.MODEL pmod pmos(vto=-1 lambda=0.02)
.MODEL nmod nmos(vto= 1 lambda=0.02)
.DC v1 0 5 0.25
.PROBE
.END