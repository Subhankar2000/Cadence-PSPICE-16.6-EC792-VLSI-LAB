123_Amrita EXP-1(a) PSPICE Three CMOS Inverters varying Kn/Kp
v1 1 0 dc 0
v2 5 0 dc 5
m1 2 1 5 5 pmod(w=10u  l=10u)
m2 3 1 5 5 pmod(w=10u  l=10u)
m3 4 1 5 5 pmod(w=10u  l=10u)
m4 2 1 0 0 nmod(w=200u l=2u)
m5 3 1 0 0 nmod(w=20u  l=2u)
m6 4 1 0 0 nmod(w=2u   l=2u)
.model pmod pmos(vto=-1 lambda=0.02)
.model nmod nmos(vto= 1 lambda=0.02)
.dc v1 0 5 0.25
.probe
.end