CMOS_INVERTER_28082020
v1 1 0 DC 0
v2 3 0 DC 5
m1 2 1 3 3 pmod(w=10u l=10u)
m2 2 1 0 0 nmod(w=10u l=10u)
.MODEL pmod pmos(vto=-1 lambda=0.02)
.MODEL nmod nmos(vto= 1 lambda=0.02)
.DC v1 0 5 0.25
.PROBE
.END